module exponentiation (
    input clk,
    input rst,
    input start,
    input [31:0] base,
    input [31:0] exponent,
    output reg [63:0] result,
    output reg done
);
    reg [7:0] count;
    reg [63:0] temp;

    always @(posedge clk or negedge rst) 
    begin
        if (!rst) 
         begin
            result <= 1;
            temp <= 0 ;
            count <= 0;
            done <= 0;
         end 
        else if (start) 
         begin
          if (count < exponent) 
             begin
                result <= result * temp;
                count <= count + 1;
             end 
           else 
              begin
                temp <= base;
                done <= 1;
            end
         end
       else
            begin
                temp <= base;
            end
    end
endmodule